library verilog;
use verilog.vl_types.all;
entity FeedForwardNN_tb is
end FeedForwardNN_tb;
